--------------------------------------------------
-- File:    decoder_scancode_ascii_tb.vhd
-- Author:  Henrique Krausburg Corrêa
--------------------------------------------------

library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all; 
    
entity decoder_scancode_ascii_tb is

	generic
	(
		CLK_EDGE    : std_logic := '1'
	);

end decoder_scancode_ascii_tb;


architecture decoder_scancode_ascii_tb of decoder_scancode_ascii_tb is

	constant	PERIOD	: time := 20 ns;										-- period time.

	-- decoder signals.
	signal 	s_scancode_in      : std_logic_vector(7 downto 0) := (others => '0');	-- scancode input (generated by input_gen)
	signal 	s_golden_ascii_out        : std_logic_vector(7 downto 0) := (others => '0');		-- decoded ascii out from golden image
	--signal 	s_cuv_ascii_out        : std_logic_vector(7 downto 0) := (others => '0');		-- decoded ascii out from cuv

begin

    --Process used to generate input values for 
	input_gen: process
	begin
		wait for PERIOD;
		s_scancode_in	<= s_scancode_in + 1;	 
	end process;

	--Instantiate golden image
	golden_decoder_scancode_ascii: entity work.decoder_scancode_ascii
	port map
	(
    	scancode_in  => s_scancode_in,		-- entrada de dados.
		ascii_out     => s_golden_ascii_out		-- Ya Yb Yc Yd Ye Yf Yg Ypto.
    );


end decoder_scancode_ascii_tb;


