--------------------------------------------------
-- File:    <nome_do_arquivo>.vhd
-- Author:  Prof. M.Sc. Marlon Moraes
-- E-mail:  marlon.moraes@pucrs.br
--------------------------------------------------


library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all; 
    
entity entity_name is

	generic
	(

	);

	port
	(
	
	);

end entity_name;


architecture architecture_name of entity_name is

    

begin



end architecture_name;


