--------------------------------------------------
-- File:    decoder_scancode_ascii_tb.vhd
-- Author:  Henrique Krausburg Corrêa
--------------------------------------------------

library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all;

library work;
    use work.txt_util.all;

entity decoder_scancode_ascii_tb is

	generic
	(
		CLK_EDGE    : std_logic := '1'
	);

end decoder_scancode_ascii_tb;


architecture decoder_scancode_ascii_tb of decoder_scancode_ascii_tb is

	constant	PERIOD	: time := 20 ns;	-- period time.
	constant	HALF_PERIOD	: time := 10 ns;	-- period time.

	-- auxiliary signals
	signal s_clk: std_logic := '1';				--Clock reference used in testbench
	signal s_finishTest: std_logic := '0';		--Flag to indicate if test finish

	-- decoder signals.
	signal 	s_scancode_in      		: std_logic_vector(7 downto 0) := (others => '0');	-- scancode input (generated by input_gen)
	signal 	s_golden_ascii_out      : std_logic_vector(7 downto 0) := (others => '0');	-- decoded ascii out from golden image
	signal 	s_cuv_ascii_out        	: std_logic_vector(7 downto 0) := (others => '0');	-- decoded ascii out from cuv

begin

	--Clock generation
	--Works untill test is not finished
	s_clk <= not s_clk after HALF_PERIOD when s_finishTest /= '1' else '0';

	--finish condition: s_scancode_in reach value x"ff"
	s_finishTest <= '1' after HALF_PERIOD when s_scancode_in = x"ff" else '0';

    --Process used to generate input values for golden and cuv blocks
	input_gen: process (s_clk)
	begin
		if(s_clk'event and s_clk = '1') then
			s_scancode_in <= s_scancode_in + 1;
		end if;
	end process;

	--Instantiate golden image
	golden_decoder_scancode_ascii: entity work.decoder_scancode_ascii
	port map
	(
    	scancode_in	=> s_scancode_in,		-- entrada de dados.
		ascii_out 	=> s_golden_ascii_out	--
    );

	--Instantiate CUV
	cuv_decoder_scancode_ascii: entity work.decoder_scancode_ascii_map
	port map
	(
    	scancode_in	=> s_scancode_in,		-- entrada de dados.
		ascii_out 	=> s_cuv_ascii_out		--
    );

	--Checker block

	checker: process (s_clk)
	begin
		if(s_clk'event and s_clk = '0') then
			assert (s_golden_ascii_out = s_cuv_ascii_out) report "CUV output is not equal to GOLDEN output. Expected: 0x" & hstr(s_golden_ascii_out) & " Got: 0x" & hstr(s_cuv_ascii_out) severity error;
		end if;
	end process;

end decoder_scancode_ascii_tb;